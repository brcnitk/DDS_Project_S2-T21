// SMART RING WITH BODY VITAL SENSORS
//S2_T21
//1. 221CS217 , Dhanush V , dhanushv.221cs217@nitk.edu.in , 9353241312
//2. 221CS222 , Harsha J Gundapalli , harshajgundapalli.221cs222@nitk.edu.in ,8792251009
//3. 221CS226 , Isiri Dinesh S , isiridineshs.221cs226@nitk.edu.in , 7349437557

module S2_T21_tb;
	reg [0:7] A; // Inputs given from the sensors
	reg [0:7] B;
	reg [0:7] C;
	reg [0:7] F1; // Fixed inputs specified in advance
	reg [0:7] F2;
	reg [0:7] F3;
	reg [0:7] F4;
	reg X;
	wire [0:7] D; // Gives us the amount of oxygen given out
	wire E; // Tells us if it is an emergency or not 
	int i;


	S2_T21 M1(A,B,C,F1,F2,F3,F4,X,D,E);


	initial 
	begin
		$dumpfile("S2_T21.vcd");
		$dumpvars(0, S2_T21_tb);
	end 

	initial
	begin 

		$display("|                S2_T21                                                                                                                               
                                                                                                   |");
		$display("----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------");
		$display("|   Input                                                                                                                                                                                                
                                        | Output-1                                              | Output-2  |");
			
	$display("-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------");
		$display("| A[0] | A[1] | A[2] | A[3] | A[4] | A[5] | A[6] | A[7] | B[0] | B[1] | B[2] | B[3] | B[4] | B[5] | B[6] | B[7] | C[0] | C[1] | C[2] | C[3] | C[4] | C[5] | C[6] | C[7] | D[0] | D[1] | D[2] | D[3] | D[4] | D[5] | D[6] | D[7] |     E     |");
		$display("-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------");
		$monitor("| %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b | %b |", A[0], A[1], A[2], A[3], A[4], A[5], A[6], A[7], B[0], B[1], B[2], B[3], B[4], B[5], B[6], B[7], C[0], C[1], C[2], C[3], C[4], C[5], C[6], C[7], D[0], D[1], D[2], D[3], D[4], D[5], D[6], D[7], E);
		

	A = 8'b00000000;
	B = 8'b00000000;
	C = 8'b00000000;
	F1 = 8'b00110111;
	F2 = 8'b01110010;
	F3 = 8'b10010101;
	F4 = 8'b00011000;
	for(i=1;i=255;i++)
	{
		#10 A = A + 8'b00000001;
		#10 B = B + 8'b00000001;
		#10 C = C + 8'b00000001;
	}
	end
	
	initial #300 $finish;


endmodule 
	
  